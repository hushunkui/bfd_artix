// Build ID Verilog Module
//
// Date:             14122019
// Time:             122541

module firmware_rev
(
   output [31:0]  firmware_date,
   output [31:0]  firmware_time
);

   assign firmware_date = 32'h14122019;
   assign firmware_time = 32'h122541;

endmodule
