// Build ID Verilog Module
//
// Date:             16122019
// Time:             213343

module firmware_rev
(
   output [31:0]  firmware_date,
   output [31:0]  firmware_time
);

   assign firmware_date = 32'h16122019;
   assign firmware_time = 32'h213343;

endmodule
