// Build ID Verilog Module
//
// Date:             09012020
// Time:             202103

module firmware_rev
(
   output [31:0]  firmware_date,
   output [31:0]  firmware_time
);

   assign firmware_date = 32'h09012020;
   assign firmware_time = 32'h202103;

endmodule
