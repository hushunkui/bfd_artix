// Build ID Verilog Module
//
// Date:             20112019
// Time:             201544

module firmware_rev
(
   output [31:0]  firmware_date,
   output [31:0]  firmware_time
);

   assign firmware_date = 32'h20112019;
   assign firmware_time = 32'h201544;

endmodule
